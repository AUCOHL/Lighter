 /*
 	Copyright 2022 AUC Open Source Hardware Lab
	
	Licensed under the Apache License, Version 2.0 (the "License"); 
	you may not use this file except in compliance with the License. 
	You may obtain a copy of the License at:

	http://www.apache.org/licenses/LICENSE-2.0

	Unless required by applicable law or agreed to in writing, software 
	distributed under the License is distributed on an "AS IS" BASIS, 
	WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
	See the License for the specific language governing permissions and 
	limitations under the License.
*/
 
 (* blackbox *)
module gf180mcu_fd_sc_mcu9t5v0__icgtp_1
    input TE,
    input E, 
    input CLK,
    output Q);
endmodule

 (* blackbox *)
module gf180mcu_fd_sc_mcu9t5v0__icgtp_2
    input TE,
    input E, 
    input CLK,
    output Q);
endmodule

 (* blackbox *)
module gf180mcu_fd_sc_mcu9t5v0__icgtp_4
    input TE,
    input E, 
    input CLK,
    output Q);
endmodule


